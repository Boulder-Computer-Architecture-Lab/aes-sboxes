/////////////////////////////////////////////////////////////////////////////////
//
// Original Author: Sumio Morioka and Akashi Satoh
// Adapted by: Phaedra Curlin
// 
// Create Date: 08/2022
// Module Name: pprm_inverter
// Project Name: aes-v
// Description: GF(2^8) inverter for the 3-Stage Positive-Polarity
//              Reed Muller S-box.
// 
// Dependencies: pprm_stage_1, pprm_stage_2, pprm_stage_3.
// 
// Revision:
// Revision 0.01 - File Created
// 
// Additional Comments: Based on design from "An Optimized S-Box Circuit
//                      Architecture for Low Power AES Design".
// 
//////////////////////////////////////////////////////////////////////////////////
`timescale 1 ns / 1 ns  // time-unit = 1 ns, precision = 1 ns

`default_nettype none

module pprm_inverter(
        input   wire    [7:0]   X,
        output  wire    [7:0]   Y
    );
    
    //----------------------------------------------------------------
    // Wires/Regs
    //----------------------------------------------------------------
    wire [3:0] A,B,C,D;

    //----------------------------------------------------------------
    // Module instantiations
    //----------------------------------------------------------------
    // PPRM Inverter Stage 1
    pprm_stage_1 stage1(
        .X(X),
        .A(A),
        .B(B),
        .C(C)
    );

    // PPRM Inverter Stage 2
    pprm_stage_2 stage2(
        .C(C),
        .D(D)
    );

    // PPRM Inverter Stage 3
    pprm_stage_3 stage3(
       .A(A),
       .B(B),
       .D(D),
       .Y(Y)
    );
    
endmodule // pprm_inverter